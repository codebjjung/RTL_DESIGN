module mcu;
endmodule

