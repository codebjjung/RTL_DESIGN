module lenet5 {
	input ap_clk,
	input ap_rst_n,
	output m_axi_memory_bus_AWVALID,
	
