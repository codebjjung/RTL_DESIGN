module pc;

